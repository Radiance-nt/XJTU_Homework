--YMQ.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY YMQ IS
  PORT(AIN4: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
       DOUT7:  OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END YMQ; 
ARCHITECTURE ART OF YMQ IS
BEGIN
  PROCESS(AIN4)
    BEGIN
    CASE AIN4 IS
    WHEN "0000"=>DOUT7<="0111111";      --0
    WHEN "0001"=>DOUT7<="0000110";      --1
    WHEN "0010"=>DOUT7<="1011011";      --2
    WHEN "0011"=>DOUT7<="1001111";      --3
    WHEN "0100"=>DOUT7<="1100110";      --4
    WHEN "0101"=>DOUT7<="1101101";      --5
    WHEN "0110"=>DOUT7<="1111101";      --6
    WHEN "0111"=>DOUT7<="0000111";      --7
    WHEN "1000"=>DOUT7<="1111111";      --8
    WHEN "1001"=>DOUT7<="1101111";      --9
    WHEN OTHERS=>DOUT7<="0000000"; 
    END CASE; 
  END PROCESS;
END ARCHITECTURE ART;